// For mode selection
`define AES256  3
`define AES196  2
`define AES128  1