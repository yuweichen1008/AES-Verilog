package aes_pkg
    `include "aes_define.sv"

    `include "aes_base.sv"
    `include "aes_encrypt.sv"
    `include "aes_decrypt.sv"

    `include "aes.sv"
endpackage